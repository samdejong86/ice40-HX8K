../common/ledscan.vhd